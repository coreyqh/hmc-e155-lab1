// TODO: fill module